comparator_inst : comparator PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		aleb	 => aleb_sig
	);
